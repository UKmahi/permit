----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:35:11 04/13/2022 
-- Design Name: 
-- Module Name:    HALFAdder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity HALFAdder is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Sum : out  STD_LOGIC;
           Carry : out  STD_LOGIC);
end HALFAdder;

architecture Behavioral of HALFAdder is

begin

 process(A,B)
  begin
  if(A ='0'and B ='0')then 
    Sum<='0';   Carry<='0';
  elsif(A ='0'and B ='1')then 
    Sum<='1'; 
	 Carry<='0';
  elsif(A ='1'and B ='0')then 
    Sum<='1'; 
	 Carry<='0';
  else   
    Sum<='0';   
	 Carry<='1';
  end if;
 end process;

end Behavioral;

